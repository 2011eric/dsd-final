module MEM(

);
endmodule